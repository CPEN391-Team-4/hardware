-- trdb_d5m.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity trdb_d5m is
	port (
		clk_sys_clk                                         : in    std_logic                     := '0';             --                                         clk_sys.clk
		clk_trdb_d5m_pixclk_clk                             : in    std_logic                     := '0';             --                             clk_trdb_d5m_pixclk.clk
		cmos_sensor_acquisition_0_cmos_sensor_input_irq_irq : out   std_logic;                                        -- cmos_sensor_acquisition_0_cmos_sensor_input_irq.irq
		i2c_scl                                             : inout std_logic                     := '0';             --                                             i2c.scl
		i2c_sda                                             : inout std_logic                     := '0';             --                                                .sda
		i2c_interrupt_sender_irq                            : out   std_logic;                                        --                            i2c_interrupt_sender.irq
		master_address                                      : out   std_logic_vector(31 downto 0);                    --                                          master.address
		master_write                                        : out   std_logic;                                        --                                                .write
		master_byteenable                                   : out   std_logic_vector(3 downto 0);                     --                                                .byteenable
		master_writedata                                    : out   std_logic_vector(31 downto 0);                    --                                                .writedata
		master_waitrequest                                  : in    std_logic                     := '0';             --                                                .waitrequest
		master_burstcount                                   : out   std_logic_vector(4 downto 0);                     --                                                .burstcount
		msgdma_csr_irq_irq                                  : out   std_logic;                                        --                                  msgdma_csr_irq.irq
		reset_reset_n                                       : in    std_logic                     := '0';             --                                           reset.reset_n
		slave_waitrequest                                   : out   std_logic;                                        --                                           slave.waitrequest
		slave_readdata                                      : out   std_logic_vector(31 downto 0);                    --                                                .readdata
		slave_readdatavalid                                 : out   std_logic;                                        --                                                .readdatavalid
		slave_burstcount                                    : in    std_logic_vector(0 downto 0)  := (others => '0'); --                                                .burstcount
		slave_writedata                                     : in    std_logic_vector(31 downto 0) := (others => '0'); --                                                .writedata
		slave_address                                       : in    std_logic_vector(6 downto 0)  := (others => '0'); --                                                .address
		slave_write                                         : in    std_logic                     := '0';             --                                                .write
		slave_read                                          : in    std_logic                     := '0';             --                                                .read
		slave_byteenable                                    : in    std_logic_vector(3 downto 0)  := (others => '0'); --                                                .byteenable
		slave_debugaccess                                   : in    std_logic                     := '0';             --                                                .debugaccess
		trdb_d5m_d_frame_valid                              : in    std_logic                     := '0';             --                                      trdb_d5m_d.frame_valid
		trdb_d5m_d_line_valid                               : in    std_logic                     := '0';             --                                                .line_valid
		trdb_d5m_d_data                                     : in    std_logic_vector(11 downto 0) := (others => '0')  --                                                .data
	);
end entity trdb_d5m;

architecture rtl of trdb_d5m is
	component trdb_d5m_cmos_sensor_acquisition_0 is
		generic (
			CMOS_SENSOR_INPUT_PIX_DEPTH      : positive := 8;
			CMOS_SENSOR_INPUT_SAMPLE_EDGE    : string   := "RISING";
			CMOS_SENSOR_INPUT_MAX_WIDTH      : positive := 1920;
			CMOS_SENSOR_INPUT_MAX_HEIGHT     : positive := 1080;
			CMOS_SENSOR_INPUT_OUTPUT_WIDTH   : positive := 32;
			CMOS_SENSOR_INPUT_FIFO_DEPTH     : positive := 32;
			CMOS_SENSOR_INPUT_DEVICE_FAMILY  : string   := "Cyclone V";
			CMOS_SENSOR_INPUT_DEBAYER_ENABLE : boolean  := false;
			CMOS_SENSOR_INPUT_PACKER_ENABLE  : boolean  := false;
			DC_FIFO_DEPTH                    : positive := 16;
			DC_FIFO_WIDTH                    : positive := 32
		);
		port (
			avalon_master_address      : out std_logic_vector(31 downto 0);                    -- address
			avalon_master_write        : out std_logic;                                        -- write
			avalon_master_byteenable   : out std_logic_vector(3 downto 0);                     -- byteenable
			avalon_master_writedata    : out std_logic_vector(31 downto 0);                    -- writedata
			avalon_master_waitrequest  : in  std_logic                     := 'X';             -- waitrequest
			avalon_master_burstcount   : out std_logic_vector(4 downto 0);                     -- burstcount
			avalon_slave_waitrequest   : out std_logic;                                        -- waitrequest
			avalon_slave_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			avalon_slave_readdatavalid : out std_logic;                                        -- readdatavalid
			avalon_slave_burstcount    : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			avalon_slave_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avalon_slave_address       : in  std_logic_vector(5 downto 0)  := (others => 'X'); -- address
			avalon_slave_write         : in  std_logic                     := 'X';             -- write
			avalon_slave_read          : in  std_logic                     := 'X';             -- read
			avalon_slave_byteenable    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			avalon_slave_debugaccess   : in  std_logic                     := 'X';             -- debugaccess
			clk_in_clk_clk             : in  std_logic                     := 'X';             -- clk
			clk_in_reset_reset_n       : in  std_logic                     := 'X';             -- reset_n
			clk_out_clk_clk            : in  std_logic                     := 'X';             -- clk
			clk_out_reset_reset_n      : in  std_logic                     := 'X';             -- reset_n
			cmos_sensor_frame_valid    : in  std_logic                     := 'X';             -- frame_valid
			cmos_sensor_line_valid     : in  std_logic                     := 'X';             -- line_valid
			cmos_sensor_data           : in  std_logic_vector(11 downto 0) := (others => 'X'); -- data
			cmos_sensor_input_irq_irq  : out std_logic;                                        -- irq
			msgdma_csr_irq_irq         : out std_logic                                         -- irq
		);
	end component trdb_d5m_cmos_sensor_acquisition_0;

	component i2c_interface is
		port (
			clk        : in    std_logic                    := 'X';             -- clk
			reset      : in    std_logic                    := 'X';             -- reset
			address    : in    std_logic_vector(1 downto 0) := (others => 'X'); -- address
			chipselect : in    std_logic                    := 'X';             -- chipselect
			write      : in    std_logic                    := 'X';             -- write
			writedata  : in    std_logic_vector(7 downto 0) := (others => 'X'); -- writedata
			read       : in    std_logic                    := 'X';             -- read
			readdata   : out   std_logic_vector(7 downto 0);                    -- readdata
			scl        : inout std_logic                    := 'X';             -- scl
			sda        : inout std_logic                    := 'X';             -- sda
			irq        : out   std_logic                                        -- irq
		);
	end component i2c_interface;

	component altera_avalon_mm_bridge is
		generic (
			DATA_WIDTH        : integer := 32;
			SYMBOL_WIDTH      : integer := 8;
			HDL_ADDR_WIDTH    : integer := 10;
			BURSTCOUNT_WIDTH  : integer := 1;
			PIPELINE_COMMAND  : integer := 1;
			PIPELINE_RESPONSE : integer := 1
		);
		port (
			clk              : in  std_logic                     := 'X';             -- clk
			reset            : in  std_logic                     := 'X';             -- reset
			s0_waitrequest   : out std_logic;                                        -- waitrequest
			s0_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			s0_readdatavalid : out std_logic;                                        -- readdatavalid
			s0_burstcount    : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			s0_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			s0_address       : in  std_logic_vector(6 downto 0)  := (others => 'X'); -- address
			s0_write         : in  std_logic                     := 'X';             -- write
			s0_read          : in  std_logic                     := 'X';             -- read
			s0_byteenable    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			s0_debugaccess   : in  std_logic                     := 'X';             -- debugaccess
			m0_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			m0_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			m0_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			m0_burstcount    : out std_logic_vector(0 downto 0);                     -- burstcount
			m0_writedata     : out std_logic_vector(31 downto 0);                    -- writedata
			m0_address       : out std_logic_vector(6 downto 0);                     -- address
			m0_write         : out std_logic;                                        -- write
			m0_read          : out std_logic;                                        -- read
			m0_byteenable    : out std_logic_vector(3 downto 0);                     -- byteenable
			m0_debugaccess   : out std_logic;                                        -- debugaccess
			s0_response      : out std_logic_vector(1 downto 0);                     -- response
			m0_response      : in  std_logic_vector(1 downto 0)  := (others => 'X')  -- response
		);
	end component altera_avalon_mm_bridge;

	component trdb_d5m_mm_interconnect_0 is
		port (
			sysclk_clk_clk                                                      : in  std_logic                     := 'X';             -- clk
			cmos_sensor_acquisition_0_clk_out_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			mm_bridge_0_reset_reset_bridge_in_reset_reset                       : in  std_logic                     := 'X';             -- reset
			mm_bridge_0_m0_address                                              : in  std_logic_vector(6 downto 0)  := (others => 'X'); -- address
			mm_bridge_0_m0_waitrequest                                          : out std_logic;                                        -- waitrequest
			mm_bridge_0_m0_burstcount                                           : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			mm_bridge_0_m0_byteenable                                           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			mm_bridge_0_m0_read                                                 : in  std_logic                     := 'X';             -- read
			mm_bridge_0_m0_readdata                                             : out std_logic_vector(31 downto 0);                    -- readdata
			mm_bridge_0_m0_readdatavalid                                        : out std_logic;                                        -- readdatavalid
			mm_bridge_0_m0_write                                                : in  std_logic                     := 'X';             -- write
			mm_bridge_0_m0_writedata                                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			mm_bridge_0_m0_debugaccess                                          : in  std_logic                     := 'X';             -- debugaccess
			cmos_sensor_acquisition_0_avalon_slave_address                      : out std_logic_vector(5 downto 0);                     -- address
			cmos_sensor_acquisition_0_avalon_slave_write                        : out std_logic;                                        -- write
			cmos_sensor_acquisition_0_avalon_slave_read                         : out std_logic;                                        -- read
			cmos_sensor_acquisition_0_avalon_slave_readdata                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			cmos_sensor_acquisition_0_avalon_slave_writedata                    : out std_logic_vector(31 downto 0);                    -- writedata
			cmos_sensor_acquisition_0_avalon_slave_burstcount                   : out std_logic_vector(0 downto 0);                     -- burstcount
			cmos_sensor_acquisition_0_avalon_slave_byteenable                   : out std_logic_vector(3 downto 0);                     -- byteenable
			cmos_sensor_acquisition_0_avalon_slave_readdatavalid                : in  std_logic                     := 'X';             -- readdatavalid
			cmos_sensor_acquisition_0_avalon_slave_waitrequest                  : in  std_logic                     := 'X';             -- waitrequest
			cmos_sensor_acquisition_0_avalon_slave_debugaccess                  : out std_logic;                                        -- debugaccess
			i2c_0_avalon_slave_address                                          : out std_logic_vector(1 downto 0);                     -- address
			i2c_0_avalon_slave_write                                            : out std_logic;                                        -- write
			i2c_0_avalon_slave_read                                             : out std_logic;                                        -- read
			i2c_0_avalon_slave_readdata                                         : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- readdata
			i2c_0_avalon_slave_writedata                                        : out std_logic_vector(7 downto 0);                     -- writedata
			i2c_0_avalon_slave_chipselect                                       : out std_logic                                         -- chipselect
		);
	end component trdb_d5m_mm_interconnect_0;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	signal mm_bridge_0_m0_waitrequest                                             : std_logic;                     -- mm_interconnect_0:mm_bridge_0_m0_waitrequest -> mm_bridge_0:m0_waitrequest
	signal mm_bridge_0_m0_readdata                                                : std_logic_vector(31 downto 0); -- mm_interconnect_0:mm_bridge_0_m0_readdata -> mm_bridge_0:m0_readdata
	signal mm_bridge_0_m0_debugaccess                                             : std_logic;                     -- mm_bridge_0:m0_debugaccess -> mm_interconnect_0:mm_bridge_0_m0_debugaccess
	signal mm_bridge_0_m0_address                                                 : std_logic_vector(6 downto 0);  -- mm_bridge_0:m0_address -> mm_interconnect_0:mm_bridge_0_m0_address
	signal mm_bridge_0_m0_read                                                    : std_logic;                     -- mm_bridge_0:m0_read -> mm_interconnect_0:mm_bridge_0_m0_read
	signal mm_bridge_0_m0_byteenable                                              : std_logic_vector(3 downto 0);  -- mm_bridge_0:m0_byteenable -> mm_interconnect_0:mm_bridge_0_m0_byteenable
	signal mm_bridge_0_m0_readdatavalid                                           : std_logic;                     -- mm_interconnect_0:mm_bridge_0_m0_readdatavalid -> mm_bridge_0:m0_readdatavalid
	signal mm_bridge_0_m0_writedata                                               : std_logic_vector(31 downto 0); -- mm_bridge_0:m0_writedata -> mm_interconnect_0:mm_bridge_0_m0_writedata
	signal mm_bridge_0_m0_write                                                   : std_logic;                     -- mm_bridge_0:m0_write -> mm_interconnect_0:mm_bridge_0_m0_write
	signal mm_bridge_0_m0_burstcount                                              : std_logic_vector(0 downto 0);  -- mm_bridge_0:m0_burstcount -> mm_interconnect_0:mm_bridge_0_m0_burstcount
	signal mm_interconnect_0_cmos_sensor_acquisition_0_avalon_slave_readdata      : std_logic_vector(31 downto 0); -- cmos_sensor_acquisition_0:avalon_slave_readdata -> mm_interconnect_0:cmos_sensor_acquisition_0_avalon_slave_readdata
	signal mm_interconnect_0_cmos_sensor_acquisition_0_avalon_slave_waitrequest   : std_logic;                     -- cmos_sensor_acquisition_0:avalon_slave_waitrequest -> mm_interconnect_0:cmos_sensor_acquisition_0_avalon_slave_waitrequest
	signal mm_interconnect_0_cmos_sensor_acquisition_0_avalon_slave_debugaccess   : std_logic;                     -- mm_interconnect_0:cmos_sensor_acquisition_0_avalon_slave_debugaccess -> cmos_sensor_acquisition_0:avalon_slave_debugaccess
	signal mm_interconnect_0_cmos_sensor_acquisition_0_avalon_slave_address       : std_logic_vector(5 downto 0);  -- mm_interconnect_0:cmos_sensor_acquisition_0_avalon_slave_address -> cmos_sensor_acquisition_0:avalon_slave_address
	signal mm_interconnect_0_cmos_sensor_acquisition_0_avalon_slave_read          : std_logic;                     -- mm_interconnect_0:cmos_sensor_acquisition_0_avalon_slave_read -> cmos_sensor_acquisition_0:avalon_slave_read
	signal mm_interconnect_0_cmos_sensor_acquisition_0_avalon_slave_byteenable    : std_logic_vector(3 downto 0);  -- mm_interconnect_0:cmos_sensor_acquisition_0_avalon_slave_byteenable -> cmos_sensor_acquisition_0:avalon_slave_byteenable
	signal mm_interconnect_0_cmos_sensor_acquisition_0_avalon_slave_readdatavalid : std_logic;                     -- cmos_sensor_acquisition_0:avalon_slave_readdatavalid -> mm_interconnect_0:cmos_sensor_acquisition_0_avalon_slave_readdatavalid
	signal mm_interconnect_0_cmos_sensor_acquisition_0_avalon_slave_write         : std_logic;                     -- mm_interconnect_0:cmos_sensor_acquisition_0_avalon_slave_write -> cmos_sensor_acquisition_0:avalon_slave_write
	signal mm_interconnect_0_cmos_sensor_acquisition_0_avalon_slave_writedata     : std_logic_vector(31 downto 0); -- mm_interconnect_0:cmos_sensor_acquisition_0_avalon_slave_writedata -> cmos_sensor_acquisition_0:avalon_slave_writedata
	signal mm_interconnect_0_cmos_sensor_acquisition_0_avalon_slave_burstcount    : std_logic_vector(0 downto 0);  -- mm_interconnect_0:cmos_sensor_acquisition_0_avalon_slave_burstcount -> cmos_sensor_acquisition_0:avalon_slave_burstcount
	signal mm_interconnect_0_i2c_0_avalon_slave_chipselect                        : std_logic;                     -- mm_interconnect_0:i2c_0_avalon_slave_chipselect -> i2c_0:chipselect
	signal mm_interconnect_0_i2c_0_avalon_slave_readdata                          : std_logic_vector(7 downto 0);  -- i2c_0:readdata -> mm_interconnect_0:i2c_0_avalon_slave_readdata
	signal mm_interconnect_0_i2c_0_avalon_slave_address                           : std_logic_vector(1 downto 0);  -- mm_interconnect_0:i2c_0_avalon_slave_address -> i2c_0:address
	signal mm_interconnect_0_i2c_0_avalon_slave_read                              : std_logic;                     -- mm_interconnect_0:i2c_0_avalon_slave_read -> i2c_0:read
	signal mm_interconnect_0_i2c_0_avalon_slave_write                             : std_logic;                     -- mm_interconnect_0:i2c_0_avalon_slave_write -> i2c_0:write
	signal mm_interconnect_0_i2c_0_avalon_slave_writedata                         : std_logic_vector(7 downto 0);  -- mm_interconnect_0:i2c_0_avalon_slave_writedata -> i2c_0:writedata
	signal rst_controller_reset_out_reset                                         : std_logic;                     -- rst_controller:reset_out -> [i2c_0:reset, mm_bridge_0:reset, mm_interconnect_0:cmos_sensor_acquisition_0_clk_out_reset_reset_bridge_in_reset_reset, mm_interconnect_0:mm_bridge_0_reset_reset_bridge_in_reset_reset]
	signal reset_reset_n_ports_inv                                                : std_logic;                     -- reset_reset_n:inv -> rst_controller:reset_in0

begin

	cmos_sensor_acquisition_0 : component trdb_d5m_cmos_sensor_acquisition_0
		generic map (
			CMOS_SENSOR_INPUT_PIX_DEPTH      => 12,
			CMOS_SENSOR_INPUT_SAMPLE_EDGE    => "FALLING",
			CMOS_SENSOR_INPUT_MAX_WIDTH      => 2592,
			CMOS_SENSOR_INPUT_MAX_HEIGHT     => 1944,
			CMOS_SENSOR_INPUT_OUTPUT_WIDTH   => 16,
			CMOS_SENSOR_INPUT_FIFO_DEPTH     => 32,
			CMOS_SENSOR_INPUT_DEVICE_FAMILY  => "Cyclone V",
			CMOS_SENSOR_INPUT_DEBAYER_ENABLE => true,
			CMOS_SENSOR_INPUT_PACKER_ENABLE  => false,
			DC_FIFO_DEPTH                    => 16,
			DC_FIFO_WIDTH                    => 32
		)
		port map (
			avalon_master_address      => master_address,                                                         --         avalon_master.address
			avalon_master_write        => master_write,                                                           --                      .write
			avalon_master_byteenable   => master_byteenable,                                                      --                      .byteenable
			avalon_master_writedata    => master_writedata,                                                       --                      .writedata
			avalon_master_waitrequest  => master_waitrequest,                                                     --                      .waitrequest
			avalon_master_burstcount   => master_burstcount,                                                      --                      .burstcount
			avalon_slave_waitrequest   => mm_interconnect_0_cmos_sensor_acquisition_0_avalon_slave_waitrequest,   --          avalon_slave.waitrequest
			avalon_slave_readdata      => mm_interconnect_0_cmos_sensor_acquisition_0_avalon_slave_readdata,      --                      .readdata
			avalon_slave_readdatavalid => mm_interconnect_0_cmos_sensor_acquisition_0_avalon_slave_readdatavalid, --                      .readdatavalid
			avalon_slave_burstcount    => mm_interconnect_0_cmos_sensor_acquisition_0_avalon_slave_burstcount,    --                      .burstcount
			avalon_slave_writedata     => mm_interconnect_0_cmos_sensor_acquisition_0_avalon_slave_writedata,     --                      .writedata
			avalon_slave_address       => mm_interconnect_0_cmos_sensor_acquisition_0_avalon_slave_address,       --                      .address
			avalon_slave_write         => mm_interconnect_0_cmos_sensor_acquisition_0_avalon_slave_write,         --                      .write
			avalon_slave_read          => mm_interconnect_0_cmos_sensor_acquisition_0_avalon_slave_read,          --                      .read
			avalon_slave_byteenable    => mm_interconnect_0_cmos_sensor_acquisition_0_avalon_slave_byteenable,    --                      .byteenable
			avalon_slave_debugaccess   => mm_interconnect_0_cmos_sensor_acquisition_0_avalon_slave_debugaccess,   --                      .debugaccess
			clk_in_clk_clk             => clk_trdb_d5m_pixclk_clk,                                                --            clk_in_clk.clk
			clk_in_reset_reset_n       => reset_reset_n,                                                          --          clk_in_reset.reset_n
			clk_out_clk_clk            => clk_sys_clk,                                                            --           clk_out_clk.clk
			clk_out_reset_reset_n      => reset_reset_n,                                                          --         clk_out_reset.reset_n
			cmos_sensor_frame_valid    => trdb_d5m_d_frame_valid,                                                 --           cmos_sensor.frame_valid
			cmos_sensor_line_valid     => trdb_d5m_d_line_valid,                                                  --                      .line_valid
			cmos_sensor_data           => trdb_d5m_d_data,                                                        --                      .data
			cmos_sensor_input_irq_irq  => cmos_sensor_acquisition_0_cmos_sensor_input_irq_irq,                    -- cmos_sensor_input_irq.irq
			msgdma_csr_irq_irq         => msgdma_csr_irq_irq                                                      --        msgdma_csr_irq.irq
		);

	i2c_0 : component i2c_interface
		port map (
			clk        => clk_sys_clk,                                     --            clock.clk
			reset      => rst_controller_reset_out_reset,                  --            reset.reset
			address    => mm_interconnect_0_i2c_0_avalon_slave_address,    --     avalon_slave.address
			chipselect => mm_interconnect_0_i2c_0_avalon_slave_chipselect, --                 .chipselect
			write      => mm_interconnect_0_i2c_0_avalon_slave_write,      --                 .write
			writedata  => mm_interconnect_0_i2c_0_avalon_slave_writedata,  --                 .writedata
			read       => mm_interconnect_0_i2c_0_avalon_slave_read,       --                 .read
			readdata   => mm_interconnect_0_i2c_0_avalon_slave_readdata,   --                 .readdata
			scl        => i2c_scl,                                         --              i2c.scl
			sda        => i2c_sda,                                         --                 .sda
			irq        => i2c_interrupt_sender_irq                         -- interrupt_sender.irq
		);

	mm_bridge_0 : component altera_avalon_mm_bridge
		generic map (
			DATA_WIDTH        => 32,
			SYMBOL_WIDTH      => 8,
			HDL_ADDR_WIDTH    => 7,
			BURSTCOUNT_WIDTH  => 1,
			PIPELINE_COMMAND  => 1,
			PIPELINE_RESPONSE => 1
		)
		port map (
			clk              => clk_sys_clk,                    --   clk.clk
			reset            => rst_controller_reset_out_reset, -- reset.reset
			s0_waitrequest   => slave_waitrequest,              --    s0.waitrequest
			s0_readdata      => slave_readdata,                 --      .readdata
			s0_readdatavalid => slave_readdatavalid,            --      .readdatavalid
			s0_burstcount    => slave_burstcount,               --      .burstcount
			s0_writedata     => slave_writedata,                --      .writedata
			s0_address       => slave_address,                  --      .address
			s0_write         => slave_write,                    --      .write
			s0_read          => slave_read,                     --      .read
			s0_byteenable    => slave_byteenable,               --      .byteenable
			s0_debugaccess   => slave_debugaccess,              --      .debugaccess
			m0_waitrequest   => mm_bridge_0_m0_waitrequest,     --    m0.waitrequest
			m0_readdata      => mm_bridge_0_m0_readdata,        --      .readdata
			m0_readdatavalid => mm_bridge_0_m0_readdatavalid,   --      .readdatavalid
			m0_burstcount    => mm_bridge_0_m0_burstcount,      --      .burstcount
			m0_writedata     => mm_bridge_0_m0_writedata,       --      .writedata
			m0_address       => mm_bridge_0_m0_address,         --      .address
			m0_write         => mm_bridge_0_m0_write,           --      .write
			m0_read          => mm_bridge_0_m0_read,            --      .read
			m0_byteenable    => mm_bridge_0_m0_byteenable,      --      .byteenable
			m0_debugaccess   => mm_bridge_0_m0_debugaccess,     --      .debugaccess
			s0_response      => open,                           -- (terminated)
			m0_response      => "00"                            -- (terminated)
		);

	mm_interconnect_0 : component trdb_d5m_mm_interconnect_0
		port map (
			sysclk_clk_clk                                                      => clk_sys_clk,                                                            --                                                    sysclk_clk.clk
			cmos_sensor_acquisition_0_clk_out_reset_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,                                         -- cmos_sensor_acquisition_0_clk_out_reset_reset_bridge_in_reset.reset
			mm_bridge_0_reset_reset_bridge_in_reset_reset                       => rst_controller_reset_out_reset,                                         --                       mm_bridge_0_reset_reset_bridge_in_reset.reset
			mm_bridge_0_m0_address                                              => mm_bridge_0_m0_address,                                                 --                                                mm_bridge_0_m0.address
			mm_bridge_0_m0_waitrequest                                          => mm_bridge_0_m0_waitrequest,                                             --                                                              .waitrequest
			mm_bridge_0_m0_burstcount                                           => mm_bridge_0_m0_burstcount,                                              --                                                              .burstcount
			mm_bridge_0_m0_byteenable                                           => mm_bridge_0_m0_byteenable,                                              --                                                              .byteenable
			mm_bridge_0_m0_read                                                 => mm_bridge_0_m0_read,                                                    --                                                              .read
			mm_bridge_0_m0_readdata                                             => mm_bridge_0_m0_readdata,                                                --                                                              .readdata
			mm_bridge_0_m0_readdatavalid                                        => mm_bridge_0_m0_readdatavalid,                                           --                                                              .readdatavalid
			mm_bridge_0_m0_write                                                => mm_bridge_0_m0_write,                                                   --                                                              .write
			mm_bridge_0_m0_writedata                                            => mm_bridge_0_m0_writedata,                                               --                                                              .writedata
			mm_bridge_0_m0_debugaccess                                          => mm_bridge_0_m0_debugaccess,                                             --                                                              .debugaccess
			cmos_sensor_acquisition_0_avalon_slave_address                      => mm_interconnect_0_cmos_sensor_acquisition_0_avalon_slave_address,       --                        cmos_sensor_acquisition_0_avalon_slave.address
			cmos_sensor_acquisition_0_avalon_slave_write                        => mm_interconnect_0_cmos_sensor_acquisition_0_avalon_slave_write,         --                                                              .write
			cmos_sensor_acquisition_0_avalon_slave_read                         => mm_interconnect_0_cmos_sensor_acquisition_0_avalon_slave_read,          --                                                              .read
			cmos_sensor_acquisition_0_avalon_slave_readdata                     => mm_interconnect_0_cmos_sensor_acquisition_0_avalon_slave_readdata,      --                                                              .readdata
			cmos_sensor_acquisition_0_avalon_slave_writedata                    => mm_interconnect_0_cmos_sensor_acquisition_0_avalon_slave_writedata,     --                                                              .writedata
			cmos_sensor_acquisition_0_avalon_slave_burstcount                   => mm_interconnect_0_cmos_sensor_acquisition_0_avalon_slave_burstcount,    --                                                              .burstcount
			cmos_sensor_acquisition_0_avalon_slave_byteenable                   => mm_interconnect_0_cmos_sensor_acquisition_0_avalon_slave_byteenable,    --                                                              .byteenable
			cmos_sensor_acquisition_0_avalon_slave_readdatavalid                => mm_interconnect_0_cmos_sensor_acquisition_0_avalon_slave_readdatavalid, --                                                              .readdatavalid
			cmos_sensor_acquisition_0_avalon_slave_waitrequest                  => mm_interconnect_0_cmos_sensor_acquisition_0_avalon_slave_waitrequest,   --                                                              .waitrequest
			cmos_sensor_acquisition_0_avalon_slave_debugaccess                  => mm_interconnect_0_cmos_sensor_acquisition_0_avalon_slave_debugaccess,   --                                                              .debugaccess
			i2c_0_avalon_slave_address                                          => mm_interconnect_0_i2c_0_avalon_slave_address,                           --                                            i2c_0_avalon_slave.address
			i2c_0_avalon_slave_write                                            => mm_interconnect_0_i2c_0_avalon_slave_write,                             --                                                              .write
			i2c_0_avalon_slave_read                                             => mm_interconnect_0_i2c_0_avalon_slave_read,                              --                                                              .read
			i2c_0_avalon_slave_readdata                                         => mm_interconnect_0_i2c_0_avalon_slave_readdata,                          --                                                              .readdata
			i2c_0_avalon_slave_writedata                                        => mm_interconnect_0_i2c_0_avalon_slave_writedata,                         --                                                              .writedata
			i2c_0_avalon_slave_chipselect                                       => mm_interconnect_0_i2c_0_avalon_slave_chipselect                         --                                                              .chipselect
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,        -- reset_in0.reset
			clk            => clk_sys_clk,                    --       clk.clk
			reset_out      => rst_controller_reset_out_reset, -- reset_out.reset
			reset_req      => open,                           -- (terminated)
			reset_req_in0  => '0',                            -- (terminated)
			reset_in1      => '0',                            -- (terminated)
			reset_req_in1  => '0',                            -- (terminated)
			reset_in2      => '0',                            -- (terminated)
			reset_req_in2  => '0',                            -- (terminated)
			reset_in3      => '0',                            -- (terminated)
			reset_req_in3  => '0',                            -- (terminated)
			reset_in4      => '0',                            -- (terminated)
			reset_req_in4  => '0',                            -- (terminated)
			reset_in5      => '0',                            -- (terminated)
			reset_req_in5  => '0',                            -- (terminated)
			reset_in6      => '0',                            -- (terminated)
			reset_req_in6  => '0',                            -- (terminated)
			reset_in7      => '0',                            -- (terminated)
			reset_req_in7  => '0',                            -- (terminated)
			reset_in8      => '0',                            -- (terminated)
			reset_req_in8  => '0',                            -- (terminated)
			reset_in9      => '0',                            -- (terminated)
			reset_req_in9  => '0',                            -- (terminated)
			reset_in10     => '0',                            -- (terminated)
			reset_req_in10 => '0',                            -- (terminated)
			reset_in11     => '0',                            -- (terminated)
			reset_req_in11 => '0',                            -- (terminated)
			reset_in12     => '0',                            -- (terminated)
			reset_req_in12 => '0',                            -- (terminated)
			reset_in13     => '0',                            -- (terminated)
			reset_req_in13 => '0',                            -- (terminated)
			reset_in14     => '0',                            -- (terminated)
			reset_req_in14 => '0',                            -- (terminated)
			reset_in15     => '0',                            -- (terminated)
			reset_req_in15 => '0'                             -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

end architecture rtl; -- of trdb_d5m
