-- system.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity system is
	port (
		clk_clk                          : in    std_logic                     := '0';             --                  clk.clk
		reset_reset_n                    : in    std_logic                     := '0';             --                reset.reset_n
		sdram_clk_clk                    : out   std_logic;                                        --            sdram_clk.clk
		sdram_controller_addr            : out   std_logic_vector(12 downto 0);                    --     sdram_controller.addr
		sdram_controller_ba              : out   std_logic_vector(1 downto 0);                     --                     .ba
		sdram_controller_cas_n           : out   std_logic;                                        --                     .cas_n
		sdram_controller_cke             : out   std_logic;                                        --                     .cke
		sdram_controller_cs_n            : out   std_logic;                                        --                     .cs_n
		sdram_controller_dq              : inout std_logic_vector(15 downto 0) := (others => '0'); --                     .dq
		sdram_controller_dqm             : out   std_logic_vector(1 downto 0);                     --                     .dqm
		sdram_controller_ras_n           : out   std_logic;                                        --                     .ras_n
		sdram_controller_we_n            : out   std_logic;                                        --                     .we_n
		trdb_d5m_cmos_sensor_frame_valid : in    std_logic                     := '0';             -- trdb_d5m_cmos_sensor.frame_valid
		trdb_d5m_cmos_sensor_line_valid  : in    std_logic                     := '0';             --                     .line_valid
		trdb_d5m_cmos_sensor_data        : in    std_logic_vector(11 downto 0) := (others => '0'); --                     .data
		trdb_d5m_i2c_scl                 : inout std_logic                     := '0';             --         trdb_d5m_i2c.scl
		trdb_d5m_i2c_sda                 : inout std_logic                     := '0';             --                     .sda
		trdb_d5m_pixclk_clk              : in    std_logic                     := '0';             --      trdb_d5m_pixclk.clk
		trdb_d5m_xclkin_clk              : out   std_logic                                         --      trdb_d5m_xclkin.clk
	);
end entity system;

architecture rtl of system is
	component system_jtag_uart_0 is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component system_jtag_uart_0;

	component system_nios2_gen2_0 is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(27 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(27 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component system_nios2_gen2_0;

	component system_pll_0 is
		port (
			refclk   : in  std_logic := 'X'; -- clk
			rst      : in  std_logic := 'X'; -- reset
			outclk_0 : out std_logic;        -- clk
			outclk_1 : out std_logic;        -- clk
			outclk_2 : out std_logic;        -- clk
			locked   : out std_logic         -- export
		);
	end component system_pll_0;

	component system_sdram_controller_0 is
		port (
			clk            : in    std_logic                     := 'X';             -- clk
			reset_n        : in    std_logic                     := 'X';             -- reset_n
			az_addr        : in    std_logic_vector(24 downto 0) := (others => 'X'); -- address
			az_be_n        : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable_n
			az_cs          : in    std_logic                     := 'X';             -- chipselect
			az_data        : in    std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			az_rd_n        : in    std_logic                     := 'X';             -- read_n
			az_wr_n        : in    std_logic                     := 'X';             -- write_n
			za_data        : out   std_logic_vector(15 downto 0);                    -- readdata
			za_valid       : out   std_logic;                                        -- readdatavalid
			za_waitrequest : out   std_logic;                                        -- waitrequest
			zs_addr        : out   std_logic_vector(12 downto 0);                    -- export
			zs_ba          : out   std_logic_vector(1 downto 0);                     -- export
			zs_cas_n       : out   std_logic;                                        -- export
			zs_cke         : out   std_logic;                                        -- export
			zs_cs_n        : out   std_logic;                                        -- export
			zs_dq          : inout std_logic_vector(15 downto 0) := (others => 'X'); -- export
			zs_dqm         : out   std_logic_vector(1 downto 0);                     -- export
			zs_ras_n       : out   std_logic;                                        -- export
			zs_we_n        : out   std_logic                                         -- export
		);
	end component system_sdram_controller_0;

	component system_trdb_d5m_0 is
		port (
			clk_sys_clk                                         : in    std_logic                     := 'X';             -- clk
			clk_trdb_d5m_pixclk_clk                             : in    std_logic                     := 'X';             -- clk
			cmos_sensor_acquisition_0_cmos_sensor_input_irq_irq : out   std_logic;                                        -- irq
			i2c_scl                                             : inout std_logic                     := 'X';             -- scl
			i2c_sda                                             : inout std_logic                     := 'X';             -- sda
			i2c_interrupt_sender_irq                            : out   std_logic;                                        -- irq
			master_address                                      : out   std_logic_vector(31 downto 0);                    -- address
			master_write                                        : out   std_logic;                                        -- write
			master_byteenable                                   : out   std_logic_vector(3 downto 0);                     -- byteenable
			master_writedata                                    : out   std_logic_vector(31 downto 0);                    -- writedata
			master_waitrequest                                  : in    std_logic                     := 'X';             -- waitrequest
			master_burstcount                                   : out   std_logic_vector(4 downto 0);                     -- burstcount
			msgdma_csr_irq_irq                                  : out   std_logic;                                        -- irq
			reset_reset_n                                       : in    std_logic                     := 'X';             -- reset_n
			slave_waitrequest                                   : out   std_logic;                                        -- waitrequest
			slave_readdata                                      : out   std_logic_vector(31 downto 0);                    -- readdata
			slave_readdatavalid                                 : out   std_logic;                                        -- readdatavalid
			slave_burstcount                                    : in    std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			slave_writedata                                     : in    std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			slave_address                                       : in    std_logic_vector(6 downto 0)  := (others => 'X'); -- address
			slave_write                                         : in    std_logic                     := 'X';             -- write
			slave_read                                          : in    std_logic                     := 'X';             -- read
			slave_byteenable                                    : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			slave_debugaccess                                   : in    std_logic                     := 'X';             -- debugaccess
			trdb_d5m_d_frame_valid                              : in    std_logic                     := 'X';             -- frame_valid
			trdb_d5m_d_line_valid                               : in    std_logic                     := 'X';             -- line_valid
			trdb_d5m_d_data                                     : in    std_logic_vector(11 downto 0) := (others => 'X')  -- data
		);
	end component system_trdb_d5m_0;

	component system_mm_interconnect_0 is
		port (
			pll_0_outclk0_clk                              : in  std_logic                     := 'X';             -- clk
			nios2_gen2_0_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			trdb_d5m_0_reset_reset_bridge_in_reset_reset   : in  std_logic                     := 'X';             -- reset
			nios2_gen2_0_data_master_address               : in  std_logic_vector(27 downto 0) := (others => 'X'); -- address
			nios2_gen2_0_data_master_waitrequest           : out std_logic;                                        -- waitrequest
			nios2_gen2_0_data_master_byteenable            : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			nios2_gen2_0_data_master_read                  : in  std_logic                     := 'X';             -- read
			nios2_gen2_0_data_master_readdata              : out std_logic_vector(31 downto 0);                    -- readdata
			nios2_gen2_0_data_master_write                 : in  std_logic                     := 'X';             -- write
			nios2_gen2_0_data_master_writedata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			nios2_gen2_0_data_master_debugaccess           : in  std_logic                     := 'X';             -- debugaccess
			nios2_gen2_0_instruction_master_address        : in  std_logic_vector(27 downto 0) := (others => 'X'); -- address
			nios2_gen2_0_instruction_master_waitrequest    : out std_logic;                                        -- waitrequest
			nios2_gen2_0_instruction_master_read           : in  std_logic                     := 'X';             -- read
			nios2_gen2_0_instruction_master_readdata       : out std_logic_vector(31 downto 0);                    -- readdata
			trdb_d5m_0_master_address                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			trdb_d5m_0_master_waitrequest                  : out std_logic;                                        -- waitrequest
			trdb_d5m_0_master_burstcount                   : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- burstcount
			trdb_d5m_0_master_byteenable                   : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			trdb_d5m_0_master_write                        : in  std_logic                     := 'X';             -- write
			trdb_d5m_0_master_writedata                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			jtag_uart_0_avalon_jtag_slave_address          : out std_logic_vector(0 downto 0);                     -- address
			jtag_uart_0_avalon_jtag_slave_write            : out std_logic;                                        -- write
			jtag_uart_0_avalon_jtag_slave_read             : out std_logic;                                        -- read
			jtag_uart_0_avalon_jtag_slave_readdata         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_uart_0_avalon_jtag_slave_writedata        : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_uart_0_avalon_jtag_slave_waitrequest      : in  std_logic                     := 'X';             -- waitrequest
			jtag_uart_0_avalon_jtag_slave_chipselect       : out std_logic;                                        -- chipselect
			nios2_gen2_0_debug_mem_slave_address           : out std_logic_vector(8 downto 0);                     -- address
			nios2_gen2_0_debug_mem_slave_write             : out std_logic;                                        -- write
			nios2_gen2_0_debug_mem_slave_read              : out std_logic;                                        -- read
			nios2_gen2_0_debug_mem_slave_readdata          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			nios2_gen2_0_debug_mem_slave_writedata         : out std_logic_vector(31 downto 0);                    -- writedata
			nios2_gen2_0_debug_mem_slave_byteenable        : out std_logic_vector(3 downto 0);                     -- byteenable
			nios2_gen2_0_debug_mem_slave_waitrequest       : in  std_logic                     := 'X';             -- waitrequest
			nios2_gen2_0_debug_mem_slave_debugaccess       : out std_logic;                                        -- debugaccess
			sdram_controller_0_s1_address                  : out std_logic_vector(24 downto 0);                    -- address
			sdram_controller_0_s1_write                    : out std_logic;                                        -- write
			sdram_controller_0_s1_read                     : out std_logic;                                        -- read
			sdram_controller_0_s1_readdata                 : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			sdram_controller_0_s1_writedata                : out std_logic_vector(15 downto 0);                    -- writedata
			sdram_controller_0_s1_byteenable               : out std_logic_vector(1 downto 0);                     -- byteenable
			sdram_controller_0_s1_readdatavalid            : in  std_logic                     := 'X';             -- readdatavalid
			sdram_controller_0_s1_waitrequest              : in  std_logic                     := 'X';             -- waitrequest
			sdram_controller_0_s1_chipselect               : out std_logic;                                        -- chipselect
			trdb_d5m_0_slave_address                       : out std_logic_vector(6 downto 0);                     -- address
			trdb_d5m_0_slave_write                         : out std_logic;                                        -- write
			trdb_d5m_0_slave_read                          : out std_logic;                                        -- read
			trdb_d5m_0_slave_readdata                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			trdb_d5m_0_slave_writedata                     : out std_logic_vector(31 downto 0);                    -- writedata
			trdb_d5m_0_slave_burstcount                    : out std_logic_vector(0 downto 0);                     -- burstcount
			trdb_d5m_0_slave_byteenable                    : out std_logic_vector(3 downto 0);                     -- byteenable
			trdb_d5m_0_slave_readdatavalid                 : in  std_logic                     := 'X';             -- readdatavalid
			trdb_d5m_0_slave_waitrequest                   : in  std_logic                     := 'X';             -- waitrequest
			trdb_d5m_0_slave_debugaccess                   : out std_logic                                         -- debugaccess
		);
	end component system_mm_interconnect_0;

	component system_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			receiver2_irq : in  std_logic                     := 'X'; -- irq
			receiver3_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component system_irq_mapper;

	component altera_irq_clock_crosser is
		generic (
			IRQ_WIDTH : integer := 1
		);
		port (
			receiver_clk   : in  std_logic                    := 'X';             -- clk
			sender_clk     : in  std_logic                    := 'X';             -- clk
			receiver_reset : in  std_logic                    := 'X';             -- reset
			sender_reset   : in  std_logic                    := 'X';             -- reset
			receiver_irq   : in  std_logic_vector(0 downto 0) := (others => 'X'); -- irq
			sender_irq     : out std_logic_vector(0 downto 0)                     -- irq
		);
	end component altera_irq_clock_crosser;

	component system_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			reset_in1      : in  std_logic := 'X'; -- reset_in1.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_req      : out std_logic;        --          .reset_req
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component system_rst_controller;

	component system_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			reset_in1      : in  std_logic := 'X'; -- reset_in1.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req      : out std_logic;
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component system_rst_controller_001;

	signal pll_0_outclk0_clk                                               : std_logic;                     -- pll_0:outclk_0 -> [irq_mapper:clk, irq_synchronizer:receiver_clk, irq_synchronizer:sender_clk, jtag_uart_0:clk, mm_interconnect_0:pll_0_outclk0_clk, nios2_gen2_0:clk, rst_controller:clk, sdram_controller_0:clk, trdb_d5m_0:clk_sys_clk]
	signal nios2_gen2_0_data_master_readdata                               : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_gen2_0_data_master_readdata -> nios2_gen2_0:d_readdata
	signal nios2_gen2_0_data_master_waitrequest                            : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_data_master_waitrequest -> nios2_gen2_0:d_waitrequest
	signal nios2_gen2_0_data_master_debugaccess                            : std_logic;                     -- nios2_gen2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_0_data_master_debugaccess
	signal nios2_gen2_0_data_master_address                                : std_logic_vector(27 downto 0); -- nios2_gen2_0:d_address -> mm_interconnect_0:nios2_gen2_0_data_master_address
	signal nios2_gen2_0_data_master_byteenable                             : std_logic_vector(3 downto 0);  -- nios2_gen2_0:d_byteenable -> mm_interconnect_0:nios2_gen2_0_data_master_byteenable
	signal nios2_gen2_0_data_master_read                                   : std_logic;                     -- nios2_gen2_0:d_read -> mm_interconnect_0:nios2_gen2_0_data_master_read
	signal nios2_gen2_0_data_master_write                                  : std_logic;                     -- nios2_gen2_0:d_write -> mm_interconnect_0:nios2_gen2_0_data_master_write
	signal nios2_gen2_0_data_master_writedata                              : std_logic_vector(31 downto 0); -- nios2_gen2_0:d_writedata -> mm_interconnect_0:nios2_gen2_0_data_master_writedata
	signal nios2_gen2_0_instruction_master_readdata                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_gen2_0_instruction_master_readdata -> nios2_gen2_0:i_readdata
	signal nios2_gen2_0_instruction_master_waitrequest                     : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_instruction_master_waitrequest -> nios2_gen2_0:i_waitrequest
	signal nios2_gen2_0_instruction_master_address                         : std_logic_vector(27 downto 0); -- nios2_gen2_0:i_address -> mm_interconnect_0:nios2_gen2_0_instruction_master_address
	signal nios2_gen2_0_instruction_master_read                            : std_logic;                     -- nios2_gen2_0:i_read -> mm_interconnect_0:nios2_gen2_0_instruction_master_read
	signal trdb_d5m_0_master_waitrequest                                   : std_logic;                     -- mm_interconnect_0:trdb_d5m_0_master_waitrequest -> trdb_d5m_0:master_waitrequest
	signal trdb_d5m_0_master_address                                       : std_logic_vector(31 downto 0); -- trdb_d5m_0:master_address -> mm_interconnect_0:trdb_d5m_0_master_address
	signal trdb_d5m_0_master_byteenable                                    : std_logic_vector(3 downto 0);  -- trdb_d5m_0:master_byteenable -> mm_interconnect_0:trdb_d5m_0_master_byteenable
	signal trdb_d5m_0_master_write                                         : std_logic;                     -- trdb_d5m_0:master_write -> mm_interconnect_0:trdb_d5m_0_master_write
	signal trdb_d5m_0_master_writedata                                     : std_logic_vector(31 downto 0); -- trdb_d5m_0:master_writedata -> mm_interconnect_0:trdb_d5m_0_master_writedata
	signal trdb_d5m_0_master_burstcount                                    : std_logic_vector(4 downto 0);  -- trdb_d5m_0:master_burstcount -> mm_interconnect_0:trdb_d5m_0_master_burstcount
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect      : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata        : std_logic_vector(31 downto 0); -- jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest     : std_logic;                     -- jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address         : std_logic_vector(0 downto 0);  -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read            : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write           : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata         : std_logic_vector(31 downto 0); -- nios2_gen2_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_readdata
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest      : std_logic;                     -- nios2_gen2_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_waitrequest
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess      : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_debugaccess -> nios2_gen2_0:debug_mem_slave_debugaccess
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address          : std_logic_vector(8 downto 0);  -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_address -> nios2_gen2_0:debug_mem_slave_address
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read             : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_read -> nios2_gen2_0:debug_mem_slave_read
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable       : std_logic_vector(3 downto 0);  -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_byteenable -> nios2_gen2_0:debug_mem_slave_byteenable
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write            : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_write -> nios2_gen2_0:debug_mem_slave_write
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata        : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_writedata -> nios2_gen2_0:debug_mem_slave_writedata
	signal mm_interconnect_0_sdram_controller_0_s1_chipselect              : std_logic;                     -- mm_interconnect_0:sdram_controller_0_s1_chipselect -> sdram_controller_0:az_cs
	signal mm_interconnect_0_sdram_controller_0_s1_readdata                : std_logic_vector(15 downto 0); -- sdram_controller_0:za_data -> mm_interconnect_0:sdram_controller_0_s1_readdata
	signal mm_interconnect_0_sdram_controller_0_s1_waitrequest             : std_logic;                     -- sdram_controller_0:za_waitrequest -> mm_interconnect_0:sdram_controller_0_s1_waitrequest
	signal mm_interconnect_0_sdram_controller_0_s1_address                 : std_logic_vector(24 downto 0); -- mm_interconnect_0:sdram_controller_0_s1_address -> sdram_controller_0:az_addr
	signal mm_interconnect_0_sdram_controller_0_s1_read                    : std_logic;                     -- mm_interconnect_0:sdram_controller_0_s1_read -> mm_interconnect_0_sdram_controller_0_s1_read:in
	signal mm_interconnect_0_sdram_controller_0_s1_byteenable              : std_logic_vector(1 downto 0);  -- mm_interconnect_0:sdram_controller_0_s1_byteenable -> mm_interconnect_0_sdram_controller_0_s1_byteenable:in
	signal mm_interconnect_0_sdram_controller_0_s1_readdatavalid           : std_logic;                     -- sdram_controller_0:za_valid -> mm_interconnect_0:sdram_controller_0_s1_readdatavalid
	signal mm_interconnect_0_sdram_controller_0_s1_write                   : std_logic;                     -- mm_interconnect_0:sdram_controller_0_s1_write -> mm_interconnect_0_sdram_controller_0_s1_write:in
	signal mm_interconnect_0_sdram_controller_0_s1_writedata               : std_logic_vector(15 downto 0); -- mm_interconnect_0:sdram_controller_0_s1_writedata -> sdram_controller_0:az_data
	signal mm_interconnect_0_trdb_d5m_0_slave_readdata                     : std_logic_vector(31 downto 0); -- trdb_d5m_0:slave_readdata -> mm_interconnect_0:trdb_d5m_0_slave_readdata
	signal mm_interconnect_0_trdb_d5m_0_slave_waitrequest                  : std_logic;                     -- trdb_d5m_0:slave_waitrequest -> mm_interconnect_0:trdb_d5m_0_slave_waitrequest
	signal mm_interconnect_0_trdb_d5m_0_slave_debugaccess                  : std_logic;                     -- mm_interconnect_0:trdb_d5m_0_slave_debugaccess -> trdb_d5m_0:slave_debugaccess
	signal mm_interconnect_0_trdb_d5m_0_slave_address                      : std_logic_vector(6 downto 0);  -- mm_interconnect_0:trdb_d5m_0_slave_address -> trdb_d5m_0:slave_address
	signal mm_interconnect_0_trdb_d5m_0_slave_read                         : std_logic;                     -- mm_interconnect_0:trdb_d5m_0_slave_read -> trdb_d5m_0:slave_read
	signal mm_interconnect_0_trdb_d5m_0_slave_byteenable                   : std_logic_vector(3 downto 0);  -- mm_interconnect_0:trdb_d5m_0_slave_byteenable -> trdb_d5m_0:slave_byteenable
	signal mm_interconnect_0_trdb_d5m_0_slave_readdatavalid                : std_logic;                     -- trdb_d5m_0:slave_readdatavalid -> mm_interconnect_0:trdb_d5m_0_slave_readdatavalid
	signal mm_interconnect_0_trdb_d5m_0_slave_write                        : std_logic;                     -- mm_interconnect_0:trdb_d5m_0_slave_write -> trdb_d5m_0:slave_write
	signal mm_interconnect_0_trdb_d5m_0_slave_writedata                    : std_logic_vector(31 downto 0); -- mm_interconnect_0:trdb_d5m_0_slave_writedata -> trdb_d5m_0:slave_writedata
	signal mm_interconnect_0_trdb_d5m_0_slave_burstcount                   : std_logic_vector(0 downto 0);  -- mm_interconnect_0:trdb_d5m_0_slave_burstcount -> trdb_d5m_0:slave_burstcount
	signal irq_mapper_receiver1_irq                                        : std_logic;                     -- trdb_d5m_0:i2c_interrupt_sender_irq -> irq_mapper:receiver1_irq
	signal irq_mapper_receiver2_irq                                        : std_logic;                     -- jtag_uart_0:av_irq -> irq_mapper:receiver2_irq
	signal irq_mapper_receiver3_irq                                        : std_logic;                     -- trdb_d5m_0:msgdma_csr_irq_irq -> irq_mapper:receiver3_irq
	signal nios2_gen2_0_irq_irq                                            : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> nios2_gen2_0:irq
	signal irq_mapper_receiver0_irq                                        : std_logic;                     -- irq_synchronizer:sender_irq -> irq_mapper:receiver0_irq
	signal irq_synchronizer_receiver_irq                                   : std_logic_vector(0 downto 0);  -- trdb_d5m_0:cmos_sensor_acquisition_0_cmos_sensor_input_irq_irq -> irq_synchronizer:receiver_irq
	signal rst_controller_reset_out_reset                                  : std_logic;                     -- rst_controller:reset_out -> [irq_mapper:reset, irq_synchronizer:receiver_reset, irq_synchronizer:sender_reset, mm_interconnect_0:nios2_gen2_0_reset_reset_bridge_in_reset_reset, mm_interconnect_0:trdb_d5m_0_reset_reset_bridge_in_reset_reset, rst_controller_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_reset_out_reset_req                              : std_logic;                     -- rst_controller:reset_req -> [nios2_gen2_0:reset_req, rst_translator:reset_req_in]
	signal nios2_gen2_0_debug_reset_request_reset                          : std_logic;                     -- nios2_gen2_0:debug_reset_request -> [rst_controller:reset_in1, rst_controller_001:reset_in1]
	signal rst_controller_001_reset_out_reset                              : std_logic;                     -- rst_controller_001:reset_out -> rst_controller_001_reset_out_reset:in
	signal reset_reset_n_ports_inv                                         : std_logic;                     -- reset_reset_n:inv -> [pll_0:rst, rst_controller:reset_in0, rst_controller_001:reset_in0]
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv  : std_logic;                     -- mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read:inv -> jtag_uart_0:av_read_n
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv : std_logic;                     -- mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write:inv -> jtag_uart_0:av_write_n
	signal mm_interconnect_0_sdram_controller_0_s1_read_ports_inv          : std_logic;                     -- mm_interconnect_0_sdram_controller_0_s1_read:inv -> sdram_controller_0:az_rd_n
	signal mm_interconnect_0_sdram_controller_0_s1_byteenable_ports_inv    : std_logic_vector(1 downto 0);  -- mm_interconnect_0_sdram_controller_0_s1_byteenable:inv -> sdram_controller_0:az_be_n
	signal mm_interconnect_0_sdram_controller_0_s1_write_ports_inv         : std_logic;                     -- mm_interconnect_0_sdram_controller_0_s1_write:inv -> sdram_controller_0:az_wr_n
	signal rst_controller_reset_out_reset_ports_inv                        : std_logic;                     -- rst_controller_reset_out_reset:inv -> [jtag_uart_0:rst_n, nios2_gen2_0:reset_n, sdram_controller_0:reset_n]
	signal rst_controller_001_reset_out_reset_ports_inv                    : std_logic;                     -- rst_controller_001_reset_out_reset:inv -> trdb_d5m_0:reset_reset_n

begin

	jtag_uart_0 : component system_jtag_uart_0
		port map (
			clk            => pll_0_outclk0_clk,                                               --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                        --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver2_irq                                         --               irq.irq
		);

	nios2_gen2_0 : component system_nios2_gen2_0
		port map (
			clk                                 => pll_0_outclk0_clk,                                          --                       clk.clk
			reset_n                             => rst_controller_reset_out_reset_ports_inv,                   --                     reset.reset_n
			reset_req                           => rst_controller_reset_out_reset_req,                         --                          .reset_req
			d_address                           => nios2_gen2_0_data_master_address,                           --               data_master.address
			d_byteenable                        => nios2_gen2_0_data_master_byteenable,                        --                          .byteenable
			d_read                              => nios2_gen2_0_data_master_read,                              --                          .read
			d_readdata                          => nios2_gen2_0_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => nios2_gen2_0_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => nios2_gen2_0_data_master_write,                             --                          .write
			d_writedata                         => nios2_gen2_0_data_master_writedata,                         --                          .writedata
			debug_mem_slave_debugaccess_to_roms => nios2_gen2_0_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => nios2_gen2_0_instruction_master_address,                    --        instruction_master.address
			i_read                              => nios2_gen2_0_instruction_master_read,                       --                          .read
			i_readdata                          => nios2_gen2_0_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => nios2_gen2_0_instruction_master_waitrequest,                --                          .waitrequest
			irq                                 => nios2_gen2_0_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => nios2_gen2_0_debug_reset_request_reset,                     --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                                        -- custom_instruction_master.readra
		);

	pll_0 : component system_pll_0
		port map (
			refclk   => clk_clk,                 --  refclk.clk
			rst      => reset_reset_n_ports_inv, --   reset.reset
			outclk_0 => pll_0_outclk0_clk,       -- outclk0.clk
			outclk_1 => sdram_clk_clk,           -- outclk1.clk
			outclk_2 => trdb_d5m_xclkin_clk,     -- outclk2.clk
			locked   => open                     -- (terminated)
		);

	sdram_controller_0 : component system_sdram_controller_0
		port map (
			clk            => pll_0_outclk0_clk,                                            --   clk.clk
			reset_n        => rst_controller_reset_out_reset_ports_inv,                     -- reset.reset_n
			az_addr        => mm_interconnect_0_sdram_controller_0_s1_address,              --    s1.address
			az_be_n        => mm_interconnect_0_sdram_controller_0_s1_byteenable_ports_inv, --      .byteenable_n
			az_cs          => mm_interconnect_0_sdram_controller_0_s1_chipselect,           --      .chipselect
			az_data        => mm_interconnect_0_sdram_controller_0_s1_writedata,            --      .writedata
			az_rd_n        => mm_interconnect_0_sdram_controller_0_s1_read_ports_inv,       --      .read_n
			az_wr_n        => mm_interconnect_0_sdram_controller_0_s1_write_ports_inv,      --      .write_n
			za_data        => mm_interconnect_0_sdram_controller_0_s1_readdata,             --      .readdata
			za_valid       => mm_interconnect_0_sdram_controller_0_s1_readdatavalid,        --      .readdatavalid
			za_waitrequest => mm_interconnect_0_sdram_controller_0_s1_waitrequest,          --      .waitrequest
			zs_addr        => sdram_controller_addr,                                        --  wire.export
			zs_ba          => sdram_controller_ba,                                          --      .export
			zs_cas_n       => sdram_controller_cas_n,                                       --      .export
			zs_cke         => sdram_controller_cke,                                         --      .export
			zs_cs_n        => sdram_controller_cs_n,                                        --      .export
			zs_dq          => sdram_controller_dq,                                          --      .export
			zs_dqm         => sdram_controller_dqm,                                         --      .export
			zs_ras_n       => sdram_controller_ras_n,                                       --      .export
			zs_we_n        => sdram_controller_we_n                                         --      .export
		);

	trdb_d5m_0 : component system_trdb_d5m_0
		port map (
			clk_sys_clk                                         => pll_0_outclk0_clk,                                --                                         clk_sys.clk
			clk_trdb_d5m_pixclk_clk                             => trdb_d5m_pixclk_clk,                              --                             clk_trdb_d5m_pixclk.clk
			cmos_sensor_acquisition_0_cmos_sensor_input_irq_irq => irq_synchronizer_receiver_irq(0),                 -- cmos_sensor_acquisition_0_cmos_sensor_input_irq.irq
			i2c_scl                                             => trdb_d5m_i2c_scl,                                 --                                             i2c.scl
			i2c_sda                                             => trdb_d5m_i2c_sda,                                 --                                                .sda
			i2c_interrupt_sender_irq                            => irq_mapper_receiver1_irq,                         --                            i2c_interrupt_sender.irq
			master_address                                      => trdb_d5m_0_master_address,                        --                                          master.address
			master_write                                        => trdb_d5m_0_master_write,                          --                                                .write
			master_byteenable                                   => trdb_d5m_0_master_byteenable,                     --                                                .byteenable
			master_writedata                                    => trdb_d5m_0_master_writedata,                      --                                                .writedata
			master_waitrequest                                  => trdb_d5m_0_master_waitrequest,                    --                                                .waitrequest
			master_burstcount                                   => trdb_d5m_0_master_burstcount,                     --                                                .burstcount
			msgdma_csr_irq_irq                                  => irq_mapper_receiver3_irq,                         --                                  msgdma_csr_irq.irq
			reset_reset_n                                       => rst_controller_001_reset_out_reset_ports_inv,     --                                           reset.reset_n
			slave_waitrequest                                   => mm_interconnect_0_trdb_d5m_0_slave_waitrequest,   --                                           slave.waitrequest
			slave_readdata                                      => mm_interconnect_0_trdb_d5m_0_slave_readdata,      --                                                .readdata
			slave_readdatavalid                                 => mm_interconnect_0_trdb_d5m_0_slave_readdatavalid, --                                                .readdatavalid
			slave_burstcount                                    => mm_interconnect_0_trdb_d5m_0_slave_burstcount,    --                                                .burstcount
			slave_writedata                                     => mm_interconnect_0_trdb_d5m_0_slave_writedata,     --                                                .writedata
			slave_address                                       => mm_interconnect_0_trdb_d5m_0_slave_address,       --                                                .address
			slave_write                                         => mm_interconnect_0_trdb_d5m_0_slave_write,         --                                                .write
			slave_read                                          => mm_interconnect_0_trdb_d5m_0_slave_read,          --                                                .read
			slave_byteenable                                    => mm_interconnect_0_trdb_d5m_0_slave_byteenable,    --                                                .byteenable
			slave_debugaccess                                   => mm_interconnect_0_trdb_d5m_0_slave_debugaccess,   --                                                .debugaccess
			trdb_d5m_d_frame_valid                              => trdb_d5m_cmos_sensor_frame_valid,                 --                                      trdb_d5m_d.frame_valid
			trdb_d5m_d_line_valid                               => trdb_d5m_cmos_sensor_line_valid,                  --                                                .line_valid
			trdb_d5m_d_data                                     => trdb_d5m_cmos_sensor_data                         --                                                .data
		);

	mm_interconnect_0 : component system_mm_interconnect_0
		port map (
			pll_0_outclk0_clk                              => pll_0_outclk0_clk,                                           --                            pll_0_outclk0.clk
			nios2_gen2_0_reset_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,                              -- nios2_gen2_0_reset_reset_bridge_in_reset.reset
			trdb_d5m_0_reset_reset_bridge_in_reset_reset   => rst_controller_reset_out_reset,                              --   trdb_d5m_0_reset_reset_bridge_in_reset.reset
			nios2_gen2_0_data_master_address               => nios2_gen2_0_data_master_address,                            --                 nios2_gen2_0_data_master.address
			nios2_gen2_0_data_master_waitrequest           => nios2_gen2_0_data_master_waitrequest,                        --                                         .waitrequest
			nios2_gen2_0_data_master_byteenable            => nios2_gen2_0_data_master_byteenable,                         --                                         .byteenable
			nios2_gen2_0_data_master_read                  => nios2_gen2_0_data_master_read,                               --                                         .read
			nios2_gen2_0_data_master_readdata              => nios2_gen2_0_data_master_readdata,                           --                                         .readdata
			nios2_gen2_0_data_master_write                 => nios2_gen2_0_data_master_write,                              --                                         .write
			nios2_gen2_0_data_master_writedata             => nios2_gen2_0_data_master_writedata,                          --                                         .writedata
			nios2_gen2_0_data_master_debugaccess           => nios2_gen2_0_data_master_debugaccess,                        --                                         .debugaccess
			nios2_gen2_0_instruction_master_address        => nios2_gen2_0_instruction_master_address,                     --          nios2_gen2_0_instruction_master.address
			nios2_gen2_0_instruction_master_waitrequest    => nios2_gen2_0_instruction_master_waitrequest,                 --                                         .waitrequest
			nios2_gen2_0_instruction_master_read           => nios2_gen2_0_instruction_master_read,                        --                                         .read
			nios2_gen2_0_instruction_master_readdata       => nios2_gen2_0_instruction_master_readdata,                    --                                         .readdata
			trdb_d5m_0_master_address                      => trdb_d5m_0_master_address,                                   --                        trdb_d5m_0_master.address
			trdb_d5m_0_master_waitrequest                  => trdb_d5m_0_master_waitrequest,                               --                                         .waitrequest
			trdb_d5m_0_master_burstcount                   => trdb_d5m_0_master_burstcount,                                --                                         .burstcount
			trdb_d5m_0_master_byteenable                   => trdb_d5m_0_master_byteenable,                                --                                         .byteenable
			trdb_d5m_0_master_write                        => trdb_d5m_0_master_write,                                     --                                         .write
			trdb_d5m_0_master_writedata                    => trdb_d5m_0_master_writedata,                                 --                                         .writedata
			jtag_uart_0_avalon_jtag_slave_address          => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address,     --            jtag_uart_0_avalon_jtag_slave.address
			jtag_uart_0_avalon_jtag_slave_write            => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write,       --                                         .write
			jtag_uart_0_avalon_jtag_slave_read             => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read,        --                                         .read
			jtag_uart_0_avalon_jtag_slave_readdata         => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata,    --                                         .readdata
			jtag_uart_0_avalon_jtag_slave_writedata        => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata,   --                                         .writedata
			jtag_uart_0_avalon_jtag_slave_waitrequest      => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest, --                                         .waitrequest
			jtag_uart_0_avalon_jtag_slave_chipselect       => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect,  --                                         .chipselect
			nios2_gen2_0_debug_mem_slave_address           => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address,      --             nios2_gen2_0_debug_mem_slave.address
			nios2_gen2_0_debug_mem_slave_write             => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write,        --                                         .write
			nios2_gen2_0_debug_mem_slave_read              => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read,         --                                         .read
			nios2_gen2_0_debug_mem_slave_readdata          => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata,     --                                         .readdata
			nios2_gen2_0_debug_mem_slave_writedata         => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata,    --                                         .writedata
			nios2_gen2_0_debug_mem_slave_byteenable        => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable,   --                                         .byteenable
			nios2_gen2_0_debug_mem_slave_waitrequest       => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest,  --                                         .waitrequest
			nios2_gen2_0_debug_mem_slave_debugaccess       => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess,  --                                         .debugaccess
			sdram_controller_0_s1_address                  => mm_interconnect_0_sdram_controller_0_s1_address,             --                    sdram_controller_0_s1.address
			sdram_controller_0_s1_write                    => mm_interconnect_0_sdram_controller_0_s1_write,               --                                         .write
			sdram_controller_0_s1_read                     => mm_interconnect_0_sdram_controller_0_s1_read,                --                                         .read
			sdram_controller_0_s1_readdata                 => mm_interconnect_0_sdram_controller_0_s1_readdata,            --                                         .readdata
			sdram_controller_0_s1_writedata                => mm_interconnect_0_sdram_controller_0_s1_writedata,           --                                         .writedata
			sdram_controller_0_s1_byteenable               => mm_interconnect_0_sdram_controller_0_s1_byteenable,          --                                         .byteenable
			sdram_controller_0_s1_readdatavalid            => mm_interconnect_0_sdram_controller_0_s1_readdatavalid,       --                                         .readdatavalid
			sdram_controller_0_s1_waitrequest              => mm_interconnect_0_sdram_controller_0_s1_waitrequest,         --                                         .waitrequest
			sdram_controller_0_s1_chipselect               => mm_interconnect_0_sdram_controller_0_s1_chipselect,          --                                         .chipselect
			trdb_d5m_0_slave_address                       => mm_interconnect_0_trdb_d5m_0_slave_address,                  --                         trdb_d5m_0_slave.address
			trdb_d5m_0_slave_write                         => mm_interconnect_0_trdb_d5m_0_slave_write,                    --                                         .write
			trdb_d5m_0_slave_read                          => mm_interconnect_0_trdb_d5m_0_slave_read,                     --                                         .read
			trdb_d5m_0_slave_readdata                      => mm_interconnect_0_trdb_d5m_0_slave_readdata,                 --                                         .readdata
			trdb_d5m_0_slave_writedata                     => mm_interconnect_0_trdb_d5m_0_slave_writedata,                --                                         .writedata
			trdb_d5m_0_slave_burstcount                    => mm_interconnect_0_trdb_d5m_0_slave_burstcount,               --                                         .burstcount
			trdb_d5m_0_slave_byteenable                    => mm_interconnect_0_trdb_d5m_0_slave_byteenable,               --                                         .byteenable
			trdb_d5m_0_slave_readdatavalid                 => mm_interconnect_0_trdb_d5m_0_slave_readdatavalid,            --                                         .readdatavalid
			trdb_d5m_0_slave_waitrequest                   => mm_interconnect_0_trdb_d5m_0_slave_waitrequest,              --                                         .waitrequest
			trdb_d5m_0_slave_debugaccess                   => mm_interconnect_0_trdb_d5m_0_slave_debugaccess               --                                         .debugaccess
		);

	irq_mapper : component system_irq_mapper
		port map (
			clk           => pll_0_outclk0_clk,              --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,       -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,       -- receiver1.irq
			receiver2_irq => irq_mapper_receiver2_irq,       -- receiver2.irq
			receiver3_irq => irq_mapper_receiver3_irq,       -- receiver3.irq
			sender_irq    => nios2_gen2_0_irq_irq            --    sender.irq
		);

	irq_synchronizer : component altera_irq_clock_crosser
		generic map (
			IRQ_WIDTH => 1
		)
		port map (
			receiver_clk   => pll_0_outclk0_clk,              --       receiver_clk.clk
			sender_clk     => pll_0_outclk0_clk,              --         sender_clk.clk
			receiver_reset => rst_controller_reset_out_reset, -- receiver_clk_reset.reset
			sender_reset   => rst_controller_reset_out_reset, --   sender_clk_reset.reset
			receiver_irq   => irq_synchronizer_receiver_irq,  --           receiver.irq
			sender_irq(0)  => irq_mapper_receiver0_irq        --             sender.irq
		);

	rst_controller : component system_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,                -- reset_in0.reset
			reset_in1      => nios2_gen2_0_debug_reset_request_reset, -- reset_in1.reset
			clk            => pll_0_outclk0_clk,                      --       clk.clk
			reset_out      => rst_controller_reset_out_reset,         -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req,     --          .reset_req
			reset_req_in0  => '0',                                    -- (terminated)
			reset_req_in1  => '0',                                    -- (terminated)
			reset_in2      => '0',                                    -- (terminated)
			reset_req_in2  => '0',                                    -- (terminated)
			reset_in3      => '0',                                    -- (terminated)
			reset_req_in3  => '0',                                    -- (terminated)
			reset_in4      => '0',                                    -- (terminated)
			reset_req_in4  => '0',                                    -- (terminated)
			reset_in5      => '0',                                    -- (terminated)
			reset_req_in5  => '0',                                    -- (terminated)
			reset_in6      => '0',                                    -- (terminated)
			reset_req_in6  => '0',                                    -- (terminated)
			reset_in7      => '0',                                    -- (terminated)
			reset_req_in7  => '0',                                    -- (terminated)
			reset_in8      => '0',                                    -- (terminated)
			reset_req_in8  => '0',                                    -- (terminated)
			reset_in9      => '0',                                    -- (terminated)
			reset_req_in9  => '0',                                    -- (terminated)
			reset_in10     => '0',                                    -- (terminated)
			reset_req_in10 => '0',                                    -- (terminated)
			reset_in11     => '0',                                    -- (terminated)
			reset_req_in11 => '0',                                    -- (terminated)
			reset_in12     => '0',                                    -- (terminated)
			reset_req_in12 => '0',                                    -- (terminated)
			reset_in13     => '0',                                    -- (terminated)
			reset_req_in13 => '0',                                    -- (terminated)
			reset_in14     => '0',                                    -- (terminated)
			reset_req_in14 => '0',                                    -- (terminated)
			reset_in15     => '0',                                    -- (terminated)
			reset_req_in15 => '0'                                     -- (terminated)
		);

	rst_controller_001 : component system_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "none",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,                -- reset_in0.reset
			reset_in1      => nios2_gen2_0_debug_reset_request_reset, -- reset_in1.reset
			clk            => open,                                   --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset,     -- reset_out.reset
			reset_req      => open,                                   -- (terminated)
			reset_req_in0  => '0',                                    -- (terminated)
			reset_req_in1  => '0',                                    -- (terminated)
			reset_in2      => '0',                                    -- (terminated)
			reset_req_in2  => '0',                                    -- (terminated)
			reset_in3      => '0',                                    -- (terminated)
			reset_req_in3  => '0',                                    -- (terminated)
			reset_in4      => '0',                                    -- (terminated)
			reset_req_in4  => '0',                                    -- (terminated)
			reset_in5      => '0',                                    -- (terminated)
			reset_req_in5  => '0',                                    -- (terminated)
			reset_in6      => '0',                                    -- (terminated)
			reset_req_in6  => '0',                                    -- (terminated)
			reset_in7      => '0',                                    -- (terminated)
			reset_req_in7  => '0',                                    -- (terminated)
			reset_in8      => '0',                                    -- (terminated)
			reset_req_in8  => '0',                                    -- (terminated)
			reset_in9      => '0',                                    -- (terminated)
			reset_req_in9  => '0',                                    -- (terminated)
			reset_in10     => '0',                                    -- (terminated)
			reset_req_in10 => '0',                                    -- (terminated)
			reset_in11     => '0',                                    -- (terminated)
			reset_req_in11 => '0',                                    -- (terminated)
			reset_in12     => '0',                                    -- (terminated)
			reset_req_in12 => '0',                                    -- (terminated)
			reset_in13     => '0',                                    -- (terminated)
			reset_req_in13 => '0',                                    -- (terminated)
			reset_in14     => '0',                                    -- (terminated)
			reset_req_in14 => '0',                                    -- (terminated)
			reset_in15     => '0',                                    -- (terminated)
			reset_req_in15 => '0'                                     -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;

	mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;

	mm_interconnect_0_sdram_controller_0_s1_read_ports_inv <= not mm_interconnect_0_sdram_controller_0_s1_read;

	mm_interconnect_0_sdram_controller_0_s1_byteenable_ports_inv <= not mm_interconnect_0_sdram_controller_0_s1_byteenable;

	mm_interconnect_0_sdram_controller_0_s1_write_ports_inv <= not mm_interconnect_0_sdram_controller_0_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

	rst_controller_001_reset_out_reset_ports_inv <= not rst_controller_001_reset_out_reset;

end architecture rtl; -- of system
